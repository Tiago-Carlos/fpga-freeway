module render (clk, cima, baixo, row, column, saida_galinha, saida_carro);
	
	input clk, cima, baixo;
	input [9:0] row, column;
	output reg saida_galinha, saida_carro;
	integer reset = 0;
	integer coluna_galinha = 320; /*column_count*/
	integer linha_galinha = 435; /*row_count*/
	
	/*tr�s carros e uma moto*/
	integer coluna_carro1 = 600;
	integer linha_carro1 = 60;
	
	integer coluna_carro2 = 0;
	integer linha_carro2 = 180;
	
	integer coluna_carro3 = 600;
	integer linha_carro3 = 300;
	
	integer coluna_moto = 600;
	integer linha_moto = 380;
	
	always @*
	begin
		/*Renderizar Galinha*/
		if(row < linha_galinha + 30 & linha_galinha < row & column < coluna_galinha + 30 & coluna_galinha < column)
			saida_galinha = 1;
		else
			saida_galinha = 0;
			
		/*Renderizar veiculos*/
		if ((row < linha_carro1 + 40 & linha_carro1 < row & column < coluna_carro1 + 60 & coluna_carro1 < column)
			|| (row < linha_carro2 + 40 & linha_carro2 < row & column < coluna_carro2 + 60 & coluna_carro2 < column)
			|| (row < linha_carro3 + 40 & linha_carro3 < row & column < coluna_carro3 + 60 & coluna_carro3 < column)
			|| (row < linha_moto + 40 & linha_moto < row & column < coluna_moto + 60 & coluna_moto < column))
			saida_carro = 1;
		else 
			saida_carro = 0;

		if ((saida_carro == 1) && (saida_galinha == 1))
			reset = 1;
	end

	// Controle for linha galinha
	always @(posedge clk)
	begin
		if(reset == 1)
			linha_galinha = 435;
		
		else if(cima == 1)
			linha_galinha = linha_galinha - 60;
			
		else if(baixo == 1)
			linha_galinha = linha_galinha + 60;
				
		if(linha_galinha >= 480) 
			linha_galinha = 435;
			
		else if(linha_galinha <= 0)
			linha_galinha = linha_galinha;
	end
	
	always @(posedge clk)
	begin
		/*Carro 1 come�a na direita da tela, e se move pra esquerda*/
		/*Velocidade 2*/
		coluna_carro1 = coluna_carro1 - 2;
		if (coluna_carro1 <= 0)
			coluna_carro1 = 640;

		/*Carro 2 come�a na esquerda da tela, e se move pra direita*/
		/*Velocidade 3*/
		coluna_carro2 = coluna_carro2 + 2;
		if (coluna_carro2 >= 640)
			coluna_carro2 = 0;

		/*Carro 3 come�a na direita da tela, e se move pra esquerda*/
		/*Velocidade 1*/
		coluna_carro3 = coluna_carro3 - 1;
		if (coluna_carro3 <= 0)
			coluna_carro3 = 640;

		/*Carro 1 come�a na direita da tela, e se move pra esquerda*/
		/*Velocidade 4*/
		coluna_moto = coluna_moto + 4;
		if (coluna_moto <= 0)
			coluna_moto = 640;
	end
	
	
	
endmodule 

/*
	4'b0011 FRENTE
	4'b1100 BAIXO
	4'b0001 TRAS
	4'b0100 CIMA
*/